/* Copyright 2020 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 * 
 * Dual Modular Redundancy Checker
 * Compares the outputs generated by two IPs and returns error signals
 * in case of mismatch
 * 
 */

module DMR_checker #(
  parameter type check_bus_t = logic,
  parameter int unsigned Pipeline  = 0,
  parameter bit AxiBus = 1'b0,
  parameter bit AxiHasAce = 1'b0
)(
  input  logic       clk_i,
  input  logic       rst_ni,
  input  check_bus_t inp_a_i,
  input  check_bus_t inp_b_i,
  output check_bus_t check_o,
  output logic       error_o
);

check_bus_t compare;
check_bus_t inp_q;
logic error;

if (AxiBus == 1) begin: gen_axi_checker
  logic error_aw, error_w, error_ar, error_r, error_b, error_ac, error_cr, error_cd;
  if (Pipeline) begin
    always_ff @(posedge clk_i, negedge rst_ni) begin
      if (~rst_ni) begin
        compare <= '0;
        inp_q   <= '0;
      end else begin
        compare.aw       <= inp_a_i.aw ^ inp_b_i.aw;
        compare.aw_valid <= inp_a_i.aw_valid ^ inp_b_i.aw_valid;
        compare.w        <= inp_a_i.w ^ inp_b_i.w;
        compare.w_valid  <= inp_a_i.w_valid ^ inp_b_i.w_valid;
        compare.ar       <= inp_a_i.ar ^ inp_b_i.ar;
        compare.ar_valid <= inp_a_i.ar_valid ^ inp_b_i.ar_valid;
        compare.r_ready  <= inp_a_i.r_ready ^ inp_b_i.r_ready;
        compare.b_ready  <= inp_a_i.b_ready ^ inp_b_i.b_ready;
        if (AxiHasAce) begin
          compare.ac_ready  <= inp_a_i.ac_ready ^ inp_b_i.ac_ready;
          compare.cr_valid  <= inp_a_i.cr_valid ^ inp_b_i.cr_valid;
          compare.cr_resp  <= inp_a_i.cr_resp ^ inp_b_i.cr_resp;
          compare.cd_valid  <= inp_a_i.cd_valid ^ inp_b_i.cd_valid;
          compare.cd  <= inp_a_i.cd ^ inp_b_i.cd;
        end
        inp_q <= inp_a_i;
      end
    end
  end else begin
    assign compare.aw       = inp_a_i.aw ^ inp_b_i.aw;
    assign compare.aw_valid = inp_a_i.aw_valid ^ inp_b_i.aw_valid;
    assign compare.w        = inp_a_i.w ^ inp_b_i.w;
    assign compare.w_valid  = inp_a_i.w_valid ^ inp_b_i.w_valid;
    assign compare.ar       = inp_a_i.ar ^ inp_b_i.ar;
    assign compare.ar_valid = inp_a_i.ar_valid ^ inp_b_i.ar_valid;
    assign compare.r_ready  = inp_a_i.r_ready ^ inp_b_i.r_ready;
    assign compare.b_ready  = inp_a_i.b_ready ^ inp_b_i.b_ready;
    if (AxiHasAce) begin
      assign compare.ac_ready  = inp_a_i.ac_ready ^ inp_b_i.ac_ready;
      assign compare.cr_valid  = inp_a_i.cr_valid ^ inp_b_i.cr_valid;
      assign compare.cr_resp  = inp_a_i.cr_resp ^ inp_b_i.cr_resp;
      assign compare.cd_valid  = inp_a_i.cd_valid ^ inp_b_i.cd_valid;
      assign compare.cd  = inp_a_i.cd ^ inp_b_i.cd;
    end
    assign inp_q = inp_a_i;
  end
  assign error_aw = (|compare.aw) | compare.aw_valid;
  assign error_w  = (|compare.w) | compare.w_valid;
  assign error_ar = (|compare.ar) | compare.ar_valid;
  assign error_r = compare.r_ready;
  assign error_b = compare.b_ready;
  if (AxiHasAce) begin
    assign error_ac  = compare.ac_ready;
    assign error_cr  = (|compare.cr_resp) | compare.cr_valid;
    assign error_cd  = (|compare.cd) | compare.cd_valid;
  end else begin
    assign error_ac  = '0;
    assign error_cr  = '0;
    assign error_cd  = '0;
  end
  assign error = error_aw | error_w | error_ar | error_r | error_b | error_ac | error_cr | error_cd;
end else begin: gen_generic_checker
  if (Pipeline) begin
    always_ff @(posedge clk_i, negedge rst_ni) begin
      if (~rst_ni) begin
        compare <= '0;
        inp_q   <= '0;
      end else begin
        compare <= inp_a_i ^ inp_b_i;
        inp_q   <= inp_a_i;
      end
    end
  end else begin
    assign compare = inp_a_i ^ inp_b_i;
    assign inp_q = inp_a_i;
  end
  assign error = |compare;
end
assign check_o = (error) ? '0 : inp_q;
assign error_o = error;

endmodule : DMR_checker
