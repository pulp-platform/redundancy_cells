// Copyright 2023 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Rapid Recovery unit with backup status registers

module rapid_recovery_unit
  import rapid_recovery_pkg::*;
#(
  parameter int unsigned RfAddrWidth     = 5,
  parameter int unsigned DataWidth       = 32,
  parameter int unsigned EccEnabled      = 1,
  parameter     type     regfile_write_t = logic,
  parameter     type     regfile_raddr_t = logic,
  parameter     type     regfile_rdata_t = logic,
  parameter     type     csr_intf_t      = logic,
  parameter     type     pc_intf_t       = logic
)(
  input  logic           clk_i,
  input  logic           rst_ni,
  /* Recovery Register File interface */
  input  regfile_write_t regfile_write_i,
  /* Recovery Control and Status Registers interface */
  input  csr_intf_t      backup_csr_i,
  output csr_intf_t      recovery_csr_o,
  /* Recovery Program Counter interface */
  input  pc_intf_t       backup_pc_i,
  output pc_intf_t       recovery_pc_o,
  /* Rapid Recovery Controller interface */
  /* backup_enable_i: result of comparison between backup_enable_o
                      (generated by the rapid_recovery_ctrl) and
                      the DMR/TMR selection mode */
  input  logic           backup_enable_i,
  /* start_recovery_i: software-requested recovery */
  input  logic           start_recovery_i,
  /* backup_enable_o: generated by rapid_recovery_ctrl, asserts that
                      the core can do the backup of its state */
  output logic           backup_enable_o,
  /* recovery_finished_o: recovery routine completion */
  output logic           recovery_finished_o,
  /* setback_o: synchronous clear for the core */
  output logic           setback_o,
  /* instr_lock_o: blocks the requests toward the instruction cache
                   during the recovery routine */
  output logic           instr_lock_o,
  /* enable_pc_recovery_o: allows the program counter to be reloaded
                           into the core */
  output logic           enable_pc_recovery_o,
  /* enable_rf_recovery_o: allows the register file to be reloaded
                           into the core */
  output logic           enable_rf_recovery_o,
  /* regfile_recovery_wdata_o: used by the address generator in the 
                               rapid_recovery_ctrl to propagate the RF
                               addresses to the core during the recovery 
                               routine */
  output regfile_write_t regfile_recovery_wdata_o, // To cores RF interface
  /* regfile_recovery_rdata_o: propagates the content from the backup RF to
                               the core RF during the recovery routine */
  output regfile_rdata_t regfile_recovery_rdata_o,
  /* debug_halt_i: signals that the cores in recovery are halted */
  input  logic           debug_halt_i,
  /* debug_req_o: sends the cores in debug mode during the recovery routine */
  output logic           debug_req_o,
  /* debug_resume_o: resumes the cores in recovery from the debug mode */
  output logic           debug_resume_o
);

logic csr_renable;

hmr_rapid_recovery_ctrl #(
  .RFAddrWidth           ( RfAddrWidth     ),
  .regfile_write_t       ( regfile_write_t )
) i_rapid_recovery_ctrl  (
  .clk_i,
  .rst_ni,
  .start_recovery_i,
  .recovery_finished_o,
  .setback_o,
  .instr_lock_o,
  .debug_req_o,
  .debug_halt_i,
  .debug_resume_o,
  .recovery_regfile_waddr_o ( regfile_recovery_wdata_o ),
  .backup_enable_o          ( backup_enable_o          ),
  .recover_csr_enable_o     ( csr_renable              ),
  .recover_pc_enable_o      ( enable_pc_recovery_o     ),
  .recover_rf_enable_o      ( enable_rf_recovery_o     )
);

recovery_csr #(
  .ECCEnabled    ( EccEnabled ),
  .csr_intf_t    ( csr_intf_t )
) i_recovery_csr (
  .clk_i,
  .rst_ni,
  .read_enable_i  ( csr_renable     ),
  .write_enable_i ( backup_enable_i ),
  .backup_csr_i   ( backup_csr_i    ),
  .recovery_csr_o ( recovery_csr_o  )
);

recovery_pc #(
  .ECCEnabled   ( EccEnabled ),
  .pc_intf_t    ( pc_intf_t  )
) i_recovery_pc (
  // Control Ports
  .clk_i,
  .rst_ni,
  .clear_i                    ( '0                   ),
  .read_enable_i              ( enable_pc_recovery_o ),
  .write_enable_i             ( backup_enable_i      ),
  // Backup Ports
  .backup_program_counter_i   ( backup_pc_i.program_counter ),
  .backup_branch_i            ( backup_pc_i.is_branch       ),
  .backup_branch_addr_i       ( backup_pc_i.branch_addr     ),
  // Recovery Pors
  .recovery_program_counter_o ( recovery_pc_o.program_counter ),
  .recovery_branch_o          ( recovery_pc_o.is_branch       ),
  .recovery_branch_addr_o     ( recovery_pc_o.branch_addr     )
);

recovery_rf  #(
  .ECCEnabled      ( EccEnabled      ),
  .ADDR_WIDTH      ( RfAddrWidth     ),
  .regfile_write_t ( regfile_write_t ),
  .regfile_raddr_t ( regfile_raddr_t ),
  .regfile_rdata_t ( regfile_rdata_t )
) i_recovery_rf    (
  .clk_i,
  .rst_ni,
  //Read port A
  .raddr_a_i    ( regfile_recovery_wdata_o.waddr_a ),
  .rdata_a_o    ( regfile_recovery_rdata_o.rdata_a ),
  //Read port B
  .raddr_b_i    ( regfile_recovery_wdata_o.waddr_b ),
  .rdata_b_o    ( regfile_recovery_rdata_o.rdata_b ),
  //Read port C
  .raddr_c_i    ( '0                                     ),
  .rdata_c_o    (                                        ),
  // Write Port A
  .waddr_a_i    ( regfile_write_i.waddr_a                ),
  .wdata_a_i    ( regfile_write_i.wdata_a                ),
  .we_a_i       ( regfile_write_i.we_a & backup_enable_i ),
  // Write Port B
  .waddr_b_i    ( regfile_write_i.waddr_b                ),
  .wdata_b_i    ( regfile_write_i.wdata_b                ),
  .we_b_i       ( regfile_write_i.we_b & backup_enable_i )
);

endmodule: rapid_recovery_unit
