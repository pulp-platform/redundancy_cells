// Copyright 2021 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Description: Testbench for the ecc register module
// Note: This testbench may only be run with the fault injection script running concurrently
// Use the 'tb_ecc_reg_multi' below to run multiple test simultaneously.

`include "ECC_reg/ecc_calc.svh"

module tb_ecc_reg #(
  parameter int unsigned DataWidth = 32,
  // ECC Settings
  parameter int unsigned NumErrorDetect = 2,
  parameter int unsigned NumErrorCorrect = 1,
  parameter bit Decode = 1,
  parameter bit Encode = 1,
  parameter bit SelfCorrect = 1,
  // FF Settings
  parameter bit HasReset = 1,
  parameter bit AsynchronousReset = 1,
  parameter bit ActiveLowReset = 1,
  parameter bit HasLoad = 0,
  // Testbench Settings
  parameter int unsigned RunCycles = 100
) (
  input  logic       enable_i,
  output logic       finished_o,
  output logic[31:0] num_errors_o
);
  // ECC dist and width calculations
  localparam int unsigned EccDist = `ECC_DIST(NumErrorCorrect, NumErrorDetect);
  localparam int          EccWidth = `ECC_WIDTH(DataWidth, EccDist);
  localparam int unsigned InputWidth  = DataWidth + (Encode ? 0 : EccWidth);
  localparam int unsigned OutputWidth = DataWidth + (Decode ? 0 : EccWidth);

  /******************
   *  Helper tasks  *
   ******************/

  localparam time         TTest     = 8ns;
  localparam time         TApply    = 2ns;

  task cycle_start();
    #TApply;
  endtask : cycle_start

  task cycle_end();
    #TTest;
  endtask : cycle_end

  /**********************
   *  Helper variables  *
   **********************/

  longint test_cnt;
  longint error_cnt;

  logic clk;
  logic rst_n;

  clk_rst_gen #(
    .ClkPeriod    ( TTest + TApply ),
    .RstClkCycles ( 5              )
  ) i_clk_gen (
    .clk_o  ( clk   ),
    .rst_no ( rst_n )
  );

  /************************
   *  Stimuli generation  *
   ************************/

  // Data type
  typedef logic [  DataWidth-1:0]        data_t;
  typedef logic [ InputWidth-1:0]        data_in_t;
  typedef logic [OutputWidth-1:0]        data_out_t;
  typedef logic [DataWidth+EccWidth-1:0] prot_t;

  class stimuli_t;
    // fixed stimuli inputs
    int num_flips;

    // randomized inputs
    rand data_t in;
    rand prot_t inject;

    constraint error_bits {$countones(inject) == num_flips;}

  endclass : stimuli_t

  // Stimuli
  stimuli_t stimuli_queue [$];

  // Golden values
  typedef struct packed {
    data_t out;
    logic e_cor, e_uncor;
  } result_t;
  result_t golden_queue[$];

  function automatic void generate_stimuli();
    // No valid output in the first cycle
    golden_queue.push_back('{out: {OutputWidth{1'b?}}, e_cor: 1'b?, e_uncor: 1'b?});

    // Step 1: No injected errors
    for (int i = 0; i < RunCycles; i++) begin
      automatic stimuli_t stimuli = new;

      stimuli.num_flips = 0;

      // Randomize
      if (!stimuli.randomize()) $error("Could not randomize.");

      stimuli_queue.push_back(stimuli);
      if(Decode) begin
        golden_queue.push_back('{out: stimuli.in, e_cor: 1'b0, e_uncor: 1'b0});
      end else begin
        golden_queue.push_back('{out: {{EccWidth{1'b?}}, stimuli.in}, e_cor: 1'b0, e_uncor: 1'b0});
      end
    end

    // Step 2: Correctable Errors
    for (int c = 1; c <= NumErrorCorrect; c++) begin
      for (int i = 0; i < RunCycles; i++) begin
        // Stimuli with fault
        automatic stimuli_t stimuli = new;
        automatic stimuli_t stimuli2 = new;
        stimuli.num_flips = c;
        if (!stimuli.randomize()) $error("Could not randomize.");

        stimuli_queue.push_back(stimuli);
        if(Decode) begin
          golden_queue.push_back('{out: stimuli.in, e_cor: 1'b1, e_uncor: 1'b0});
        end else begin
          if(stimuli.inject[DataWidth-1:0] == 0) begin
            golden_queue.push_back('{out: {{EccWidth{1'b?}}, stimuli.in}, e_cor: 1'b1, e_uncor: 1'b0});
          end else begin
            golden_queue.push_back('{out: {OutputWidth{1'b?}}, e_cor: 1'b1, e_uncor: 1'b0});
          end
        end

        // For self-correction enabled: Second stimuli without fault while error is corrected
        stimuli2.num_flips = 0;
        if (!stimuli2.randomize()) $error("Could not randomize.");

        stimuli_queue.push_back(stimuli2);
        if(Decode) begin
          if(SelfCorrect) begin
            golden_queue.push_back('{out: stimuli.in, e_cor: 1'b0, e_uncor: 1'b0});
          end else begin
            golden_queue.push_back('{out: stimuli2.in, e_cor: 1'b0, e_uncor: 1'b0});
          end
        end else begin
          if(SelfCorrect) begin
            golden_queue.push_back('{out: {{EccWidth{1'b?}}, stimuli.in}, e_cor: 1'b0, e_uncor: 1'b0});
          end else begin
            golden_queue.push_back('{out: {OutputWidth{1'b?}}, e_cor: 1'b0, e_uncor: 1'b0});
          end
        end
      end
    end

    // Step 3: Uncorrectable, Detectable Errors
    for (int c = NumErrorCorrect + 1; c <= NumErrorDetect; c++) begin
      for (int i = 0; i < RunCycles; i++) begin
        // Stimuli with fault
        automatic stimuli_t stimuli = new;
        stimuli.num_flips = c;
        if (!stimuli.randomize()) $error("Could not randomize.");

        stimuli_queue.push_back(stimuli);
        golden_queue.push_back('{out: {OutputWidth{1'b?}}, e_cor: 1'b0, e_uncor: 1'b1});
      end
    end
  endfunction : generate_stimuli

  // Apply stimuli
  data_in_t in;
  data_t in_uncoded;
  prot_t fault_mask_next, fault_mask, inject_val;

  task automatic apply_stimuli();
    automatic stimuli_t stimuli;

    wait (stimuli_queue.size() != '0);

    stimuli = stimuli_queue.pop_front();
    in_uncoded = stimuli.in;
    fault_mask_next = stimuli.inject;
  endtask : apply_stimuli

  initial begin : init_stimuli
    in_uncoded = '0;
    fault_mask_next = '0;
  end : init_stimuli

  if(!Encode) begin
    ecc_enc #(
      .DataWidth       (DataWidth      ),
      .NumErrorDetect  (NumErrorDetect ),
      .NumErrorCorrect (NumErrorCorrect)
    ) i_enc (
      .data_i (in_uncoded),
      .data_o (in        )
    );
  end else begin
    assign in = in_uncoded;
  end

  /***********************
   *  Device Under Test  *
   ***********************/

  data_out_t out;
  logic e_cor, e_uncor;

  ecc_reg #(
    .DataWidth         (DataWidth),
    .NumErrorDetect    (NumErrorDetect),
    .NumErrorCorrect   (NumErrorCorrect),
    .Encode            (Encode),
    .Decode            (Decode),
    .SelfCorrect       (SelfCorrect),
    .HasReset          (HasReset),
    .AsynchronousReset (AsynchronousReset),
    .ActiveLowReset    (ActiveLowReset),
    .HasLoad           (HasLoad)
  ) i_dut (
    .clk_i                 (clk),
    .rst_ni                (rst_n),
    .data_i                (in),
    .data_o                (out),
    .error_correctable_o   (e_cor),
    .error_uncorrectable_o (e_uncor),
    .load_en_i             ('0)
  );

  always_ff @( posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      fault_mask <= '0;
    end else begin
      fault_mask <= fault_mask_next;
    end
  end

  assign inject_val = fault_mask ^ i_dut.data_q;

  /***********************
   *  Output collection  *
   ***********************/

  result_t result_queue [$];

  function automatic void collect_result;
    result_queue.push_back('{out: out,e_cor: e_cor, e_uncor: e_uncor});
  endfunction: collect_result

  task automatic check_result;
    automatic result_t result;
    automatic result_t golden;

    do begin
      wait(result_queue.size() != 0);

      // Capture the results
      result = result_queue.pop_front();
      golden = golden_queue.pop_front();

      // Account for this check
      test_cnt++;

      if (result != golden) begin
        $warning("ERROR! Test %0d: expected %p, found %p.", test_cnt, golden, result);
        error_cnt++;
      end
    end while (stimuli_queue.size() != 0);
  endtask: check_result

  /****************
   *  Test bench  *
   ****************/

  task run();
    // Apply stimuli and collect results cycle
    forever begin
      if(enable_i) begin
        cycle_start();
        apply_stimuli();
        cycle_end();
        collect_result();
      end
    end
  endtask : run

  assign num_errors_o = error_cnt;

  initial begin: tb
    // Initialize variables
    test_cnt  = '0;
    error_cnt = '0;
    finished_o = '0;

    wait(enable_i);

    $display("Generating Stimuli for Datawidth %d", DataWidth);

    @(posedge rst_n)

    fork
      // Run the TB
      run();
      fork
        // Generate stimuli
        generate_stimuli();
        // Check result
        check_result();
      join
    join_any

    finished_o = 1'b1;
  end: tb

endmodule

module tb_ecc_reg_multi #(
  parameter int unsigned MaxDataWidth = 0,
  // ECC Settings
  parameter int unsigned NumErrorDetect = 2,
  parameter int unsigned NumErrorCorrect = 1,
  parameter bit Decode = 1,
  parameter bit Encode = 1,
  parameter bit SelfCorrect = 1,
  // FF Settings
  parameter bit HasReset = 1,
  parameter bit AsynchronousReset = 1,
  parameter bit ActiveLowReset = 1,
  parameter bit HasLoad = 0,
  // Testbench parameters
  parameter int unsigned RunCycles = 50
);

  logic                         enable;
  logic[MaxDataWidth-1:0]       finished;
  logic[MaxDataWidth-1:0][31:0] error_cnt;

  for(genvar datawidth = 1; datawidth <= MaxDataWidth; datawidth++) begin : gen_dut
    tb_ecc_reg #(
      .DataWidth         (datawidth        ),
      .NumErrorDetect    (NumErrorDetect   ),
      .NumErrorCorrect   (NumErrorCorrect  ),
      .Decode            (Decode           ),
      .Encode            (Encode           ),
      .SelfCorrect       (SelfCorrect      ),
      .HasReset          (HasReset         ),
      .AsynchronousReset (AsynchronousReset),
      .ActiveLowReset    (ActiveLowReset   ),
      .HasLoad           (HasLoad          ),
      .RunCycles         (RunCycles        )
    ) i_dut (
      .enable_i     (enable                ),
      .finished_o   (finished[datawidth-1] ),
      .num_errors_o (error_cnt[datawidth-1])
    );
  end

  longint total_errors;

  initial begin
    $display("Testing With Parameters:");
    $display(" - MaxDataWidth:      %30d", MaxDataWidth);
    $display(" - NumErrorDetect:    %30d", NumErrorDetect);
    $display(" - NumErrorCorrect:   %30d", NumErrorCorrect);
    $display(" - Decode:            %30d", Decode);
    $display(" - Encode:            %30d", Encode);
    $display(" - SelfCorrect:       %30d", SelfCorrect);
    $display(" - HasReset:          %30d", HasReset);
    $display(" - AsynchronousReset: %30d", AsynchronousReset);
    $display(" - ActiveLowReset:    %30d", ActiveLowReset);
    $display(" - HasLoad:           %30d", HasLoad);

    enable = 1'b1;

    wait( finished == {MaxDataWidth{1'b1}} );

    total_errors = '0;

    $display("Testing Completed:");
    for(int i = 0; i < MaxDataWidth; i++) begin
      $display("Datawidth %d: %d Errors.", i+1, error_cnt[i]);
      total_errors += error_cnt[i];
    end

    $display("Finished Running %d tests over %d DataWidths", MaxDataWidth * RunCycles, MaxDataWidth);
    $display("Errors: %d", total_errors);

    $finish(0);

  end

endmodule
